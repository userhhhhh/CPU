// `include "config.v"
`include "/home/hqs123/class_code/CPU/src/config.v"
module RS_chooser(
    input wire clk,
    input wire rst,
    input wire rdy

    

);
    

endmodule