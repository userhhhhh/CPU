`include "config.v"
module cache(
    input wire clk,
    input wire rst,
    input wire rdy,

    
);
endmodule