`include "config.v"
module RS_chooser(
    input wire clk,
    input wire rst,
    input wire rdy,

    

);
    

endmodule